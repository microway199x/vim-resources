/////////////////////////////////////////////////////////// 
/// author : Micro
/// initial version :  #0.01 as first version 
/// initial date :  
/// modify engineer :
/// modify date : 
/// filename : 
/// function describe : 
/// 
////////////////////////////////////////////////////////////


module <Module-name> (
///{auto-port-define-begin
/*AUTOINOUT*/

/*AUTOINPUT*/

/*AUTOOUTPUT*/

///}auto-port-define-end

);

///{user-variable-define-begin

///}user-variable-define-end

///{auto-variable-define-begin

/*AUTOWIRE*/

/*AUTOREG*/

///}auto-variable-define-end

////////////////////////////////////////////////////////////



endmodule 

//Local Variables:
//verilog-library-flags:("-y incdir1/ -y incdir2/")
//verilog-library-directories:("." "dir1" "dir2" )
//eval: (defun upperx (name)
//          (uppercase name))
//eval: (defun tieoff (dir)
//          (if (string-equal dir "input")
//              (concat "{" vl-width "{1'b0}}")
//              ""))
//val:(setq verilog-auto-output-ignore-regexp (concat
//  "^\\("
//  "signal1_.*"
//  "\\|signal2_.*"
//  "\\)$"
//  )))
//End:

////////////////////////////////////////////////////////////
/// modify log :
/// modify engineer : modify date: version: what modified
///
////////////////////////////////////////////////////////////


